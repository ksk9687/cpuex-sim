000000000000000000000000000000000000,
010011000000000000000000000000000000,
000000000000001111110010000000000000,
000101001111111111111111110000000000,
000101001111111111101111110000000000,
000101001111101111101111100000000000,
000101001111101111101111100000000000,
000011000000001111000000000100001001,
110000000000000000000000000100001000,
000000000000000000010000000000000000,
000000000000000000100000000000000000,
000000000000000000110000000000000001,
110010010000010000000010100100010010,
000101000000101111010000110000000000,
000100000000110000100000000000000000,
000100001111010000110000000000000000,
000001000000010000010000000000000001,
110000000000000000000000000100001100,
011100000000100000000000000000000000,
110000000000000000000000000100010011,
