000000000000000000000000000000000000,
010011000000000000000000000000000000,
000000000000001111110010000000000000,
000101001111111111111111110000000000,
000101001111111111101111110000000000,
000101001111101111101111100000000000,
000101001111101111101111100000000000,
000011000000001111000000000100001001,
110000000000000000000000000100001000,
000000000000000000010000000000001010,
000011000000001111000000000100001101,
011100000000010000000000000000000000,
110000000000000000000000000100001100,
110011000000010000000000010100011011,
000010001111101111100000000000000011,
010010001111100000001111000000000000,
010010001111100000000000010000000001,
000010000000010000010000000000000001,
000011000000001111000000000100001101,
010010001111100000000000010000000010,
010000001111100000010000000000000001,
000010000000010000010000000000000010,
000011000000001111000000000100001101,
010000001111101111010000000000000010,
000101000000010000011111010000000000,
010000001111101111000000000000000000,
000001001111101111100000000000000011,
110110001111000000000000000000000000,
